library verilog;
use verilog.vl_types.all;
entity baud_test_vlg_vec_tst is
end baud_test_vlg_vec_tst;
