library verilog;
use verilog.vl_types.all;
entity projectDraft_vlg_vec_tst is
end projectDraft_vlg_vec_tst;
