library verilog;
use verilog.vl_types.all;
entity tx2_vlg_vec_tst is
end tx2_vlg_vec_tst;
