library verilog;
use verilog.vl_types.all;
entity testing_bus_vlg_vec_tst is
end testing_bus_vlg_vec_tst;
