library verilog;
use verilog.vl_types.all;
entity Tasinda_vlg_vec_tst is
end Tasinda_vlg_vec_tst;
