library verilog;
use verilog.vl_types.all;
entity testing_counter is
    port(
        pin_name1       : out    vl_logic
    );
end testing_counter;
