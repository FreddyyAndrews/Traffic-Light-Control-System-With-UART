library verilog;
use verilog.vl_types.all;
entity Tx_vlg_vec_tst is
end Tx_vlg_vec_tst;
